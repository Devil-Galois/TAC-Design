** Profile: "SCHEMATIC1-sim_layer1"  [ C:\Users\15062\Desktop\design\layer1-PSpiceFiles\SCHEMATIC1\sim_layer1.sim ] 

** Creating circuit file "sim_layer1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Cadence\Spb_data\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000n 0 
.OPTIONS ADVCONV
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
